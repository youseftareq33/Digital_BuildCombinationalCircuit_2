module pAnd(x, y, z);
input x,y;
output  z;


and and_gate(z,x,y);


endmodule